library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Convertidor is
	GENERIC(
		NBITS  : integer :=  24; -- Cantidad de bits del n�mero binario.
		NSALIDA: integer := 28  -- Cantidad de bits de salida en formato BCD.
	);
	PORT(
		num_bin: in  STD_LOGIC_VECTOR(NBITS-1   downto 0);
		num_bcd: inout STD_LOGIC_VECTOR(27 downto 0)
	);
end Convertidor;

architecture arq_Convertidor of Convertidor is
signal num :  STD_LOGIC_VECTOR(27 downto 0);
begin
	proceso_bcd: process(num_bin)
		variable z: STD_LOGIC_VECTOR(NBITS+NSALIDA-1 downto 0);
	begin
		-- Inicializaci�n de datos en cero.
		z := (others => '0');
		-- Se realizan los primeros tres corrimientos.
		z(NBITS+2 downto 3) := num_bin;
		-- Ciclo para las iteraciones restantes.
		for i in 0 to NBITS-4 loop
			-- Unidades (4 bits).
			if z(NBITS+3 downto NBITS) > 4 then
				z(NBITS+3 downto NBITS) := z(NBITS+3 downto NBITS) + 3;
			end if;
			-- Decenas (4 bits).
			if z(NBITS+7 downto NBITS+4) > 4 then
				z(NBITS+7 downto NBITS+4) := z(NBITS+7 downto NBITS+4) + 3;
			end if;
			-- Centenas (3 bits).
			if z(NBITS+11 downto NBITS+8) > 4 then
				z(NBITS+11 downto NBITS+8) := z(NBITS+11 downto NBITS+8) + 3;
			end if;				
					-- MIL (3 bits).
			if z(NBITS+15 downto NBITS+12) > 4 then
				z(NBITS+15 downto NBITS+12) := z(NBITS+15 downto NBITS+12) + 3;
			end if;
					-- DIEZ MIL (3 bits).

			if z(NBITS+19 downto NBITS+16) > 4 then
				z(NBITS+19 downto NBITS+16) := z(NBITS+19 downto NBITS+16) + 3;
			end if;
					-- CIEN MIL (3 bits).

			if z(NBITS+23 downto NBITS+20) > 4 then
				z(NBITS+23 downto NBITS+20) := z(NBITS+23 downto NBITS+20) + 3;
			end if;
					-- MILLON (3 bits).

			if z(NBITS+27 downto NBITS+24) > 4 then
				z(NBITS+27 downto NBITS+24) := z(NBITS+27 downto NBITS+24) + 3;
			end if;
			-- Corrimiento a la izquierda.
			z(NBITS+NSALIDA-1 downto 1) := z(NBITS+NSALIDA-2 downto 0);
		end loop;
		-- Pasando datos de variable Z, correspondiente a BCD.
		num <= z(NBITS+NSALIDA-1 downto NBITS);
	end process;
	process (num)
	begin 
	
	if (  num < "0000010000100000000000000000") then 
		    num_bcd<= "0000001000000000000000000000";
		elsif  (num >= "0000010000100000000000000000" and num < "0000010001000000000000000000") then 
		    num_bcd <= "0000001000010000000000000000";
		elsif (num >=  "0000010001000000000000000000" and num < "0000010001100000000000000000") then 
		    num_bcd <= "0000001000100000000000000000";
		elsif (num >=  "0000010001100000000000000000" and num < "0000010010000000000000000000") then 
		    num_bcd <= "0000001000110000000000000000";
		elsif (num >=  "0000010010000000000000000000" and num < "0000010100000000000000000000") then 
		    num_bcd <= "0000001001000000000000000000";
		elsif (num >=  "0000010100000000000000000000" and num < "0000010100100000000000000000") then
		   num_bcd <= "0000001001010000000000000000";
		elsif (num >=  "0000010100100000000000000000" and num < "0000010101000000000000000000") then
          num_bcd <= "0000001001100000000000000000";		
		elsif (num >=  "0000010101000000000000000000" and num < "0000010101100000000000000000") then
         num_bcd <= "0000001001110000000000000000";		
		elsif (num >=  "0000010101100000000000000000" and num < "0000010110000000000000000000") then
          num_bcd <= "0000001010000000000000000000";		
		elsif (num >=  "0000010110000000000000000000" and num < "0000011000000000000000000000") then
			 num_bcd <= "0000001010010000000000000000";
		elsif (num >=  "0000011000000000000000000000" and num < "0000011000100000000000000000") then
			 num_bcd <= "0000001100000000000000000000";
		elsif (num >=  "0000011000100000000000000000" and num < "0000011001000000000000000000") then
		    num_bcd <= "0000001100010000000000000000";
		elsif (num >=  "0000011001000000000000000000" and num < "0000011010000000000000000000") then
         num_bcd <= "0000001100100000000000000000";		
		elsif (num >=  "0000011010000000000000000000" and num < "0000011100000000000000000000") then
			 num_bcd <= "0000001100110000000000000000";
      elsif (num >=  "0000011100000000000000000000" and num < "0000011100100000000000000000") then
		    num_bcd <= "0000001101000000000000000000";
      elsif (num >=  "0000011100100000000000000000" and num < "0000011101000000000000000000") then
			 num_bcd <= "0000001101010000000000000000";
      elsif (num >=  "0000011101000000000000000000" and num < "0000011101100000000000000000") then
			 num_bcd <= "0000001101100000000000000000";
		elsif (num >=  "0000011101100000000000000000" and num < "0000011110000000000000000000") then
			 num_bcd <= "0000001101110000000000000000";
		elsif (num >=  "0000011110000000000000000000" and num < "0000100000000000000000000000") then
			num_bcd <= "0000001110000000000000000000";
		elsif (num >=  "0000100000000000000000000000" and num < "0000100000100000000000000000") then
		    num_bcd <= "0000001110010000000000000000";
		elsif (num >=  "0000100000100000000000000000" and num < "0000100001000000000000000000") then 
		    num_bcd <= "0000010000010000000000000000";
		elsif (num >=  "0000100001000000000000000000" and num < "0000100001100000000000000000") then
		    num_bcd <= "0000010000100000000000000000";
		elsif (num >=  "0000100001100000000000000000" and num < "0000100010000000000000000000") then 
			 num_bcd <= "0000010000110000000000000000";
		elsif (num >=  "0000100010000000000000000000" and num < "0000100100000000000000000000") then 
		    num_bcd <= "0000010001000000000000000000";
		elsif (num >=  "0000100100000000000000000000" and num < "0000100100100000000000000000") then
			 num_bcd <= "0000010001010000000000000000";
		elsif (num >=  "0000100100100000000000000000" and num < "0000100101000000000000000000") then
			 num_bcd <= "0000010001100000000000000000";
		elsif (num >=  "0000100101000000000000000000" and num < "0000100101100000000000000000") then 
		    num_bcd <= "0000010001110000000000000000";
		elsif (num >=  "0000100101100000000000000000" and num < "0000100110000000000000000000") then 
		    num_bcd <= "0000010010000000000000000000";
		elsif (num >=  "0000100110000000000000000000" and num < "0001000000000000000000000000") then
          num_bcd <= "0000010010010000000000000000";		
		elsif (num >=  "0001000000000000000000000000" and num < "0001000000100000000000000000") then 
		    num_bcd <= "0000010100000000000000000000";
		elsif (num >=  "0001000000100000000000000000" and num < "0001000001000000000000000000") then
			 num_bcd <= "0000010100010000000000000000";
		elsif (num >=  "0001000001000000000000000000" and num < "0001000001100000000000000000") then 
		    num_bcd <= "0000010100100000000000000000";
		elsif (num >=  "0001000001100000000000000000" and num < "0001000010000000000000000000") then
          num_bcd <= "0000010100110000000000000000";		
		elsif (num >=  "0001000010000000000000000000" and num < "0001000100000000000000000000") then
		    num_bcd <= "0000010101000000000000000000";
		elsif (num >=  "0001000100000000000000000000" and num < "0001000100100000000000000000") then 
		    num_bcd <= "0000010101010000000000000000";
		elsif (num >=  "0001000100100000000000000000" and num < "0001000101000000000000000000") then 
		    num_bcd <= "0000010101100000000000000000";
		elsif (num >=  "0001000101000000000000000000" and num < "0001000101100000000000000000") then 
		    num_bcd <= "0000010101110000000000000000";
		elsif (num >=  "0001000101100000000000000000" and num < "0001000110000000000000000000") then
		    num_bcd <= "0000010110000000000000000000";
		elsif (num >=  "0001000110000000000000000000" and num < "0001001000000000000000000000") then
          num_bcd <= "0000010110010000000000000000";		
		elsif (num >=  "0001001000000000000000000000" and num < "0001001000100000000000000000") then 
		    num_bcd <= "0000011000000000000000000000";
		elsif (num >=  "0001001000100000000000000000" and num < "0001001001000000000000000000") then
          num_bcd <= "0000011000010000000000000000";		
		elsif (num >=  "0001001001000000000000000000" and num < "0001001001100000000000000000") then
		    num_bcd <= "0000011000100000000000000000";
		elsif (num >=  "0001001001100000000000000000" and num < "0001001010000000000000000000") then 
		    num_bcd <= "0000011000110000000000000000";
		elsif (num >=  "0001001010000000000000000000" and num < "0001001100000000000000000000") then
		    num_bcd <= "0000011001000000000000000000";
		elsif (num >=  "0001001100000000000000000000" and num < "0001001100100000000000000000") then
		    num_bcd <= "0000011001010000000000000000";
		elsif (num >=  "0001001100100000000000000000" and num < "0001001101000000000000000000") then 
		    num_bcd <= "0000011001100000000000000000";
		elsif (num >=  "0001001101000000000000000000" and num < "0001001101100000000000000000") then
          num_bcd <= "0000011001110000000000000000";		
		elsif (num >=  "0001001101100000000000000000" and num < "0001001110000000000000000000") then
          num_bcd <= "0000011010000000000000000000";		
		elsif (num >=  "0001001110000000000000000000" and num < "0001010000000000000000000000") then
          num_bcd <= "0000011010010000000000000000";		
		elsif (num >=  "0001010000000000000000000000" and num < "0001010000100000000000000000") then 
		    num_bcd <= "0000011100000000000000000000";
		elsif (num >=  "0001010000100000000000000000" and num < "0001010001000000000000000000") then
          num_bcd <= "0000011100010000000000000000";		
		elsif (num >=  "0001010001000000000000000000" and num < "0001010001100000000000000000") then
          num_bcd <= "0000011100100000000000000000";		
	   elsif (num >=  "0001010001100000000000000000" and num < "0001010010000000000000000000") then
          num_bcd <= "0000011100110000000000000000";		
		elsif (num >=  "0001010010000000000000000000" and num < "0001010100000000000000000000") then
          num_bcd <= "0000011101000000000000000000";		
		elsif (num >=  "0001010100000000000000000000" and num < "0001010100100000000000000000") then
		    num_bcd <= "0000011101010000000000000000";
		elsif (num >=  "0001010100100000000000000000" and num < "0001010101000000000000000000") then
          num_bcd <= "0000011101100000000000000000";		
		elsif (num >=  "0001010101000000000000000000" and num < "0001010101100000000000000000") then
          num_bcd <= "0000011101110000000000000000";		
		elsif (num >=  "0001010101100000000000000000" and num < "0001010110000000000000000000") then
          num_bcd <= "0000011110000000000000000000";		
		elsif (num >=  "0001010110000000000000000000" and num < "0001011000000000000000000000") then
          num_bcd <= "0000011110010000000000000000";		
		elsif (num >=  "0001011000000000000000000000" and num < "0001011000100000000000000000") then
		    num_bcd <= "0000100000000000000000000000";
		elsif (num >=  "0001011000100000000000000000" and num < "0001011001000000000000000000") then
		    num_bcd <= "0000100000010000000000000000";
		elsif (num >=  "0001011001000000000000000000" and num < "0001011010000000000000000000") then 
		    num_bcd <= "0000100000100000000000000000";
		elsif (num >=  "0001011010000000000000000000" and num < "0001011100000000000000000000") then
	       num_bcd <= "0000100000110000000000000000";
      elsif (num >=  "0001011100000000000000000000" and num < "0001011100100000000000000000") then
	       num_bcd <= "0000100001000000000000000000";
      elsif (num >=  "0001011100100000000000000000" and num < "0001011101000000000000000000") then
          num_bcd <= "0000100001010000000000000000";		
      elsif (num >=  "0001011101000000000000000000" and num < "0001011101100000000000000000") then
          num_bcd <= "0000100001100000000000000000";		
		elsif (num >=  "0001011101100000000000000000" and num < "0001011110000000000000000000") then 
		    num_bcd <= "0000100001110000000000000000";
		elsif (num >=  "0001011110000000000000000000" and num < "0001100000000000000000000000") then
		    num_bcd <= "0000100010000000000000000000";
		elsif (num >=  "0001100000000000000000000000" and num < "0001100000100000000000000000") then
          num_bcd <= "0000100010010000000000000000";
		elsif (num >=  "0001100000100000000000000000" and num < "0001100001000000000000000000") then
          num_bcd <= "0000100100000000000000000000";		
		elsif (num >=  "0001100001000000000000000000" and num < "0001100001100000000000000000") then
		    num_bcd <= "0000100100010000000000000000";
		elsif (num >=  "0001100001100000000000000000" and num < "0001100010000000000000000000") then
          num_bcd <= "0000100100100000000000000000";		
		elsif (num >=  "0001100010000000000000000000" and num < "0001100100000000000000000000") then
          num_bcd <= "0000100100110000000000000000";		
		elsif (num >=  "0001100100000000000000000000" and num < "0001100100100000000000000000") then 
		    num_bcd <= "0000100101000000000000000000";
		elsif (num >=  "0001100100100000000000000000" and num < "0001100101000000000000000000") then
          num_bcd <= "0000100101010000000000000000";		
		elsif (num >=  "0001100101000000000000000000" and num < "0001100101100000000000000000") then
          num_bcd <= "0000100101100000000000000000";		
		elsif (num >=  "0001100101100000000000000000" and num < "0001100110000000000000000000") then 
		    num_bcd <= "0000100101110000000000000000";
		elsif (num >=  "0001100110000000000000000000" and num < "0010000000000000000000000000") then 
		    num_bcd <= "0000100110000000000000000000";
		elsif (num >=  "0010000000000000000000000000" and num < "0010000000100000000000000000") then
		    num_bcd <= "0000100110010000000000000000";
		elsif (num >=  "0010000000100000000000000000" and num < "0010000001000000000000000000") then 
	       num_bcd <= "0001000000000000000000000000";
		elsif (num >=  "0010000001000000000000000000" and num < "0010000001100000000000000000") then 
		    num_bcd <= "0001000000010000000000000000";
		elsif (num >=  "0010000001100000000000000000" and num < "0010000010000000000000000000") then
          num_bcd <= "0001000000100000000000000000";		
		elsif (num >=  "0010000010000000000000000000" and num < "0010000100000000000000000000") then 
		    num_bcd <= "0001000000110000000000000000";
		elsif (num >=  "0010000100000000000000000000" and num < "0010000100100000000000000000") then 
		    num_bcd <= "0001000001000000000000000000";
		elsif (num >=  "0010000100100000000000000000" and num < "0010000101000000000000000000") then 
		    num_bcd <= "0001000001010000000000000000";
		elsif (num >=  "0010000101000000000000000000" and num < "0010000101100000000000000000") then 
		    num_bcd <= "0001000001100000000000000000";
		elsif (num >=  "0010000101100000000000000000" and num < "0010000110000000000000000000") then
          num_bcd <= "0001000001110000000000000000";		
		elsif (num >=  "0010000110000000000000000000" and num < "0010001000000000000000000000") then 
		    num_bcd <= "0001000010010000000000000000";
		elsif (num >=  "0010001000000000000000000000" and num < "0010001000100000000000000000") then 
		    num_bcd <= "0001000100000000000000000000";
		elsif (num >=  "0010001000100000000000000000" and num < "0010001001000000000000000000") then 
		    num_bcd <= "0001000100010000000000000000";
		elsif (num >=  "0010001001000000000000000000" and num < "0010001001100000000000000000") then
		    num_bcd <= "0001000100100000000000000000";
		elsif (num >=  "0010001001100000000000000000" and num < "0010001010000000000000000000") then 
		    num_bcd <= "0001000100110000000000000000";
		elsif (num >=  "0010001010000000000000000000" and num < "0010001100000000000000000000") then
	       num_bcd <= "0001000101000000000000000000";				 
		elsif (num >=  "0010001100000000000000000000" and num < "0010001100100000000000000000") then
		    num_bcd <= "0001000101010000000000000000";
		elsif (num >=  "0010001100100000000000000000" and num < "0010001101000000000000000000") then 
	       num_bcd <= "0001000101100000000000000000";	
		elsif (num >=  "0010001101000000000000000000" and num < "0010001101100000000000000000") then 
          num_bcd <= "0001000101110000000000000000";		
		elsif (num >=  "0010001101100000000000000000" and num < "0010001110000000000000000000") then 
		    num_bcd <= "0001000110000000000000000000";
		elsif (num >=  "0010001110000000000000000000" and num < "0010010000000000000000000000") then 
		    num_bcd <= "0001000110010000000000000000";
		elsif (num >=  "0010010000000000000000000000" and num < "0010010000100000000000000000") then 
		    num_bcd <= "0001001000000000000000000000";
		elsif (num >=  "0010010000100000000000000000" and num < "0010010001000000000000000000") then 
          num_bcd <= "0001001000010000000000000000";		
		elsif (num >=  "0010010001000000000000000000" and num < "0010010001100000000000000000") then 
		    num_bcd <= "0001001000100000000000000000";
		elsif (num >=  "0010010001100000000000000000" and num < "0010010010000000000000000000") then 
		    num_bcd <= "0001001000110000000000000000";
		elsif (num >=  "0010010010000000000000000000" and num < "0010010100000000000000000000") then 
          num_bcd <= "0001001001000000000000000000";		
		elsif (num >=  "0010010100000000000000000000" and num < "0010010100100000000000000000") then
		    num_bcd <= "0001001010010000000000000000";
		elsif (num >=  "0010010100100000000000000000" and num < "0010010101000000000000000000") then 
		    num_bcd <= "0001001001100000000000000000";
		elsif (num >=  "0010010101000000000000000000" and num < "0010010101100000000000000000") then 
          num_bcd <= "0001001001110000000000000000";		
		elsif (num >=  "0010010101100000000000000000" and num < "0010010110000000000000000000") then 
		    num_bcd <= "0001001010000000000000000000";
		elsif (num >=  "0010010110000000000000000000" and num < "0010011000000000000000000000") then 
		    num_bcd <= "0001001010010000000000000000";
		elsif (num >=  "0010011000000000000000000000" and num < "0010011000100000000000000000") then 
		    num_bcd <= "0001001100000000000000000000";
		elsif (num >=  "0010011000100000000000000000" and num < "0010011001000000000000000000") then
          num_bcd <= "0001001100010000000000000000";		
		elsif (num >=  "0010011001000000000000000000" and num < "0010011010000000000000000000") then 
		    num_bcd <= "0001001100100000000000000000";
		elsif (num >=  "0010011010000000000000000000" and num < "0010011100000000000000000000") then
          num_bcd <= "0001001100110000000000000000";
		elsif (num >=  "0010011100000000000000000000" and num < "0010011100100000000000000000") then
          num_bcd <= "0001001101000000000000000000";
		elsif (num >=  "0010011100100000000000000000" and num < "0010011101000000000000000000") then 
          num_bcd <= "0001001110010000000000000000";
		elsif (num >=  "0010011101000000000000000000" and num < "0010011101100000000000000000") then 
		    num_bcd <= "0001001101100000000000000000";
		elsif (num >=  "0010011101100000000000000000" and num < "0010011110000000000000000000") then 
		    num_bcd <= "0001001101110000000000000000";
		elsif (num >=  "0010011110000000000000000000" and num < "0010100000000000000000000000") then
		    num_bcd <= "0001001110000000000000000000";
		elsif (num >=  "0010100000000000000000000000" and num < "0010100000100000000000000000") then
		    num_bcd <= "0001001110010000000000000000";
		elsif (num >=  "0010100000100000000000000000" and num < "0010100001000000000000000000") then 
		    num_bcd <= "0001010000000000000000000000";
		elsif (num >=  "0010100001000000000000000000" and num < "0010100001100000000000000000") then
		    num_bcd <= "0001010000010000000000000000";
		elsif (num >=  "0010100001100000000000000000" and num < "0010100010000000000000000000") then 
		    num_bcd <= "0001010000100000000000000000";
		elsif (num >=  "0010100010000000000000000000" and num < "0010100100000000000000000000") then 
		    num_bcd <= "0001010000110000000000000000";
		elsif (num >=  "0010100100000000000000000000") then
		    num_bcd <= "0001010001000000000000000000";
		else
		num_bcd <= num;
		end if;
		end process;
end arq_Convertidor;


