`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
//////////////////////////////////////////////////////////////////////////////////
module comp_sum(a,b,s);
input [7:0]a,b;//numero mayor de 255, numero mayor de 510
output


endmodule
