`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
//////////////////////////////////////////////////////////////////////////////////
module suma(a,b,s);
input [7:0]a,b;//numero mayor de 255, numero mayor de 510
output [8:0]s;//porque la suma es mas grande de 511

assign s=a+b;

endmodule
