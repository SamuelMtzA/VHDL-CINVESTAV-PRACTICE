`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
//////////////////////////////////////////////////////////////////////////////////
module sumador(a,b,cin,cout,s);
input [31:0]a,b;
input cin;
output [31:0]s;
output cout;

	assign {cout,s}=a+b+cin;//concatenar las salidas

endmodule
